driver logic
i have modified driver
