monitor logic
