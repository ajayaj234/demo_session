driver logic
