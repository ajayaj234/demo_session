generetor logic
